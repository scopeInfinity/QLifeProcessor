// `include "emulator/chipset.v"

module chipset_test;
    // wire reset; // reset button
    // CHIPSET dut(.reset(reset));

    // initial begin
    //     assign reset = 0; // button is never pressed.
    // end
endmodule
