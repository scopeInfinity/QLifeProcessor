module ADD_4_16b(
    output[15:0] out,
    input[15:0] in);

    assign out = in + 4;
endmodule
