// `include "emulator/module/mblock/mconst.v"

module MCONST_test;
//     reg[31:0] in;
//     wire[31:0] out;

//     MCONST dut(.out(out),
//         .in(in));

//     initial begin
//         in = 16'b0010111100010010;
//         # 10
//         $display("MCONST_TEST: in=%b out=%b", in, out);
//         if (out !== 32'b00000000000000000010111100010010) begin
//             $error("mconst failed");
//             $fatal(1);
//         end
//         in = 16'b1001011000011000;
//         # 10
//         $display("MCONST_TEST: in=%b out=%b", in, out);
//         if (out !== 32'b00000000000000001001011000011000) begin
//             $error("mconst failed");
//             $fatal(1);
//         end
//     end
endmodule
