module BOOT_CONTROL(output is_powered_on);
    // TODO: Needs improvement.
    assign is_powered_on = 1;
endmodule