// module ROM_boot(address, value)

// endmodule;
