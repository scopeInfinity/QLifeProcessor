`include "emulator/rom.v"

module rom_test;
reg a,b,c,d;
output e;

// ROM r(a,b,c,d,e);

// initial begin
//   a=1'b0;
//   b=1'b0;
//   d=1'b0;
//   c=1'b1;
// //   e=1'b1;
//   # 10
//   $display("a=%b b=%b c=%b d=%b e=%b", a,b,c,d,e);
//   # 10 c=1'b0;
//   # 10
//   $display("a=%b b=%b c=%b d=%b e=%b", a,b,c,d,e);
//   $monitor("a=%b b=%b c=%b d=%b e=%b", a,b,c,d,e);
//   # 10000
//   $finish;
// end

endmodule