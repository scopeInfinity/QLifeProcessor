`include "emulator/module/stag0_ins_resolver.v"
`include "emulator/module/stage1or2_store.v"

module PROCESSOR(
    output[15:0] mblock_address,
    output[31:0] mblock_input,
    output[1:0] mblock_selector,
    input[31:0] mblock_output,

    );


endmodule;
